module ram_single(
output reg [7:0] q,
input [9:0] a,
input [7:0] d,
input we, clk
);
reg [7:0] mem [1024:0];
always @(posedge clk) begin
if (we) mem[a] <= d;
q <= mem[a];
end
endmodule

module address_interface(input [9:0] in_addr, input[2:0] oper, input clk,  output [9:0] out_addr);

reg [9:0] address = 10'b0;
reg written;

always @(posedge clk)
begin
	if (oper[0] & ~written) address <= address + 10'b1;
	else if (oper[1] & ~written) address <= address - 10'b1;
	else if (oper[2] & ~written) address <= in_addr;
	else address <= address;
	written <= |oper ;
end

assign out_addr = address;

endmodule

module hex_to_seg(input [3:0] hex, output [6:0] seg);
	function [6:0] convert(input [3:0] code);
		case(code)
			4'h0: convert = 7'b1000000;
			4'h1: convert = 7'b1111001;
			4'h2: convert = 7'b0100100;
			4'h3: convert = 7'b0110000;
			4'h4: convert = 7'b0011001;
			4'h5: convert = 7'b0010010;
			4'h6: convert = 7'b0000010;
			4'h7: convert = 7'b1111000;
			4'h8: convert = 7'b0000000;
			4'h9: convert = 7'b0010000;
			4'ha: convert = 7'b0001000;
			4'hb: convert = 7'b0000011;
			4'hc: convert = 7'b1000110;
			4'hd: convert = 7'b0100001;
			4'he: convert = 7'b0000110;
			4'hf: convert = 7'b0001110;
		endcase
	endfunction

	assign seg = convert(hex);
endmodule

//=======================================================
//  This code is generated by Terasic System Builder
//=======================================================

module Memory(

	//////////// CLOCK //////////
	input 		          		CLOCK2_50,
	input 		          		CLOCK3_50,
	input 		          		CLOCK4_50,
	input 		          		CLOCK_50,

	//////////// SEG7 //////////
	output		     [6:0]		HEX0,
	output		     [6:0]		HEX1,
	output		     [6:0]		HEX2,
	output		     [6:0]		HEX3,
	output		     [6:0]		HEX4,
	output		     [6:0]		HEX5,

	//////////// KEY //////////
	input 		     [3:0]		KEY,

	//////////// LED //////////
	output		     [9:0]		LEDR,

	//////////// SW //////////
	input 		     [9:0]		SW
);



//=======================================================
//  REG/WIRE declarations
//=======================================================

wire [9:0] addr_out;
wire [7:0] data_out;
wire [2:0] oper;
reg block_write;

//=======================================================
//  Structural coding
//=======================================================

assign LEDR[7:0] = data_out;
assign LEDR[9] = addr_out[9];
assign LEDR[8] = addr_out[8];
assign oper = ~KEY[2:0];

always @(posedge CLOCK_50)
begin 
	block_write <= ~KEY[3] ? 1'b1 : 1'b0;
end

address_interface i1(.in_addr(SW[9:0]), .oper(oper), .clk(CLOCK_50), .out_addr(addr_out));
ram_single rs1(.q(data_out), .a(addr_out), .d(SW[7:0]), .we(~KEY[3] & ~block_write), .clk(CLOCK_50));

hex_to_seg addr_low(.hex(addr_out[3:0]), .seg(HEX0));
hex_to_seg addr_high(.hex(addr_out[7:4]), .seg(HEX1));

hex_to_seg data_low(.hex(data_out[3:0]), .seg(HEX2));
hex_to_seg data_high(.hex(data_out[7:4]), .seg(HEX3));

hex_to_seg sw_low(.hex(SW[3:0]), .seg(HEX4));
hex_to_seg sw_high(.hex(SW[7:4]), .seg(HEX5));

endmodule
